Checkout this file!
